module tmr_rtc #
(
  parameter FREQ = 100000000
)
(
  //----------------------------------------------------------------------------------------------------------------------
  // Inputs
  //----------------------------------------------------------------------------------------------------------------------
  input                   tmr_clk,
  input                   tmr_resetn,
  //----------------------------------------------------------------------------------------------------------------------
  // Outputs
  //----------------------------------------------------------------------------------------------------------------------
  output     [31:0]       tmr_rtc_data_out
);
  //----------------------------------------------------------------------------------------------------------------------
  // Includes
  //----------------------------------------------------------------------------------------------------------------------
  `include "tmr_func.v"

  //----------------------------------------------------------------------------------------------------------------------
  // Local Parameters
  //----------------------------------------------------------------------------------------------------------------------
  localparam [31:0] PRESC_MAX_VAL = 0.001*FREQ-1;
  localparam [31:0] PRESC_W       = log2(PRESC_MAX_VAL);
  
  //----------------------------------------------------------------------------------------------------------------------
  // Internal Signals
  //----------------------------------------------------------------------------------------------------------------------

  // Prescaler
  reg [PRESC_W-1:0] presc_reg;
  reg [31:0]        rtc_reg;

  // Real-Time CLock
  wire              rtc_en;

  //----------------------------------------------------------------------------------------------------------------------
  // Prescaler
  //----------------------------------------------------------------------------------------------------------------------
  always @ (posedge tmr_clk or negedge tmr_resetn)
    if (~tmr_resetn)
      presc_reg <= {PRESC_W{1'b0}};
    else if (presc_reg == PRESC_MAX_VAL[31:0])
      presc_reg <= {PRESC_W{1'b0}};
    else
      presc_reg <= presc_reg + {{PRESC_W-1{1'b0}}, 1'b1};
      
  assign rtc_en = presc_reg == PRESC_MAX_VAL;
  
  //----------------------------------------------------------------------------------------------------------------------
  // Real-Time Clock
  //----------------------------------------------------------------------------------------------------------------------
  always @ (posedge tmr_clk or negedge tmr_resetn)
    if (~tmr_resetn)
      rtc_reg <= 32'd0;
    else if (rtc_en)
      rtc_reg <= rtc_reg + 32'd1;
    else
      rtc_reg <= rtc_reg;
      
  assign tmr_rtc_data_out = rtc_reg;

endmodule